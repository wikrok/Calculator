----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:23:47 05/01/2017 
-- Design Name: 
-- Module Name:    DeIntegernator - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DeIntegernator is
	port(integerIn : IN INTEGER;
		  integerValid : IN STD_LOGIC;
		  enable : IN STD_LOGIC;
		  reset : IN STD_LOGIC;
		  charOut : OUT STD_LOGIC_VECTOR (7 downto 0)
		  
		  );
		  
		  

end DeIntegernator;

architecture Behavioral of DeIntegernator is

begin


end Behavioral;

